module RS2_Data_Execute_Mux (input logic [31:0] rs2_data_ex, input logic [31:0] data_to_write, input logic [31:0] address_to_write_into,
output logic [31:0] src_BE
);
